`timescale 1ns / 1ps

module tb_multiplier_top;

    localparam int PRECISION        = 8;
    localparam int BIAS_PRECISION   = 32;
    localparam int NUM_FEATURES     = 2;
    localparam int MUL_PER_FEATURE  = 16;
    localparam int N                = 16;
    localparam int M_MUL            = 16;
    localparam int Z_WEIGHTS        = 16;

    logic                        clk;
    logic                        rst;
    logic                        ce;
    logic [BIAS_PRECISION-1:0]   bias;
    logic [PRECISION-1:0]        weights_in [N-1:0];
    logic [PRECISION-1:0]        features   [NUM_FEATURES-1:0][N-1:0];
    logic [PRECISION-1:0]        out        [NUM_FEATURES-1:0];

    multiplier_top #(
        .PRECISION               ( PRECISION      ),
        .BIAS_PRECISION          ( BIAS_PRECISION ),
        .OUTPUT_STAGE_PRECISION  ( 64             ),
        .NUM_FEATURES            ( NUM_FEATURES   ),
        .MUL_PER_FEATURE         ( 8              ),
        .N                       ( N              ),
        .M_MUL                   ( 2094967296     ),
        .Z_WEIGHTS               ( 5              )
    ) dut (
        .clk                     ( clk            ),
        .rst                     ( rst            ),
        .ce                      ( ce             ),
        .bias                    ( bias           ),
        .weights_in              ( weights_in     ),
        .features                ( features       ),
        .out                     ( out            )
    );

    always #5 clk = ~clk;

    initial begin
        clk        = 0;
        rst        = 1;
        ce         = 0;
        bias       = 32'd10;
        
        weights_in <= '{default:0};
        features   <= '{default:0};

        @(posedge clk);
        rst <= 0;
        ce  <= 1;

        @(posedge clk);
        
        weights_in <= '{8'h01, 8'h02, 8'h03, 8'h04, 8'h05, 8'h06, 8'h07, 8'h08, 8'h01, 8'h02, 8'h03, 8'h04, 8'h05, 8'h06, 8'h07, 8'h08};
        
        features <= '{
            '{8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01},
            '{8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02}
        };
        
        @(posedge clk);
        
        weights_in <= '{8'h10, 8'h20, 8'h30, 8'h40, 8'h50, 8'h60, 8'h70, 8'h80, 8'h90, 8'hA0, 8'hB0, 8'hC0, 8'hD0, 8'hE0, 8'hF0, 8'h01};        
        
        features <= '{
            '{8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05, 8'h05},
            '{8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A, 8'h0A}
        };
        
        @(posedge clk);
    end

endmodule